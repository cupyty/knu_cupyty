module bin2seg(
input	wire	[3:0]	bin,

output	reg		[7:0]	seg
);

always @(bin)
begin
	case(bin)
		////////////////////////////////////////////
		4'd0 : seg = 8'b00000011
		4'd1 : seg = 8'b10011111
		4'd2 : seg = 8'b00100101
		4'd3 : seg = 8'b00001101
		4'd4 : seg = 8'b10011001
		4'd5 : seg = 8'b01001001
		4'd6 : seg = 8'b01000001
		4'd7 : seg = 8'b00011011
		4'd8 : seg = 8'b00000001
		4'd9 : seg = 8'b00011001
		4'd10 : seg = 8'b11111101
		default : seg = 8'b11111111
		////////////////////////////////////////////
	endcase
end

endmodule
